module write_byte(input wire [63:0] address,
                  input wire [7:0] data,
    
                  output reg [7:0] result);

address[]
